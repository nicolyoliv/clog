library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Declaração da entidade: Subtrator de 4 bits
entity subtractor_4bits is
    port(
        num1, num2 : in std_logic_vector(3 downto 0); -- Entradas de 4 bits
        num3 : out std_logic_vector(4 downto 0)      -- Saída de 5 bits (4 da diferença + 1 do borrow)
    );
end subtractor_4bits;

-- Arquitetura: Instancia 4 subtratores de 1 bit.
architecture subtractor_arch of subtractor_4bits is
    signal bo0, bo1, bo2, bo3 : std_logic; -- Sinais de borrow intermediários
    signal res : std_logic_vector(4 downto 0);  -- Sinal interno para o resultado
begin
    -- Subtrator do LSB (bit 0)
    subtractor_a: entity work.subtractor_1bit(subtractor_arch)
    port map(
        a => num1(0),
        b => num2(0),
        bi => '0',        -- O borrow inicial é 0
        bo => bo0,
        s => res(0)
    );
    
    -- Subtrator do bit 1, usando o borrow out do anterior
    subtractor_b: entity work.subtractor_1bit(subtractor_arch)
    port map(
        a => num1(1),
        b => num2(1),
        bi => bo0,
        bo => bo1,
        s => res(1)
        );
        
    -- Subtrator do bit 2
    subtractor_c: entity work.subtractor_1bit(subtractor_arch)
    port map(
        a => num1(2),
        b => num2(2),
        bi => bo1,
        bo => bo2,
        s => res(2)
    );
    
    -- Subtrator do MSB (bit 3)
    subtractor_d: entity work.subtractor_1bit(subtractor_arch)
    port map(
        a => num1(3),
        b => num2(3),
        bi => bo2,
        bo => res(4),   -- O borrow out final é o 5º bit do resultado
        s => res(3)
    );
    -- Atribui o resultado final, com uma lógica de underflow simplista
    num3 <= res when res(4) = '0' else
            "10000";  

end subtractor_arch;
